*scale (5), circuit type (ladderrc)

RC ladder --scale=5
VIN 1 0 1
R0 0 1 100
C0 1 0 1p
R1 1 2 100
C1 2 0 1p
R2 2 3 100
C2 3 0 1p
R3 3 4 100
C3 4 0 1p
R4 4 5 100
C4 5 0 1p
R5 5 6 100
C5 6 0 1p

.OP
.PRINT V(6)
.ends
