*scale(1)	circuit type(Clock RC tree (random fanout))

VIN 1 0 1
R0 1 2 100
C0 2 0 1p
R1 2 3 100
C1 3 0 1p
R2 3 4 100
C2 4 0 1p
R3 4 5 100
C3 5 0 1p
R4 5 6 100
C4 6 0 1p
R5 6 7 100
C5 7 0 1p
.OP
.ENDS
