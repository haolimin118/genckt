*scale(1)	circuit type(Clock R tree (random fanout))

VIN 1 0 1
R0 1 2 100
R1 2 3 100
R2 3 4 100
R3 4 5 100
R4 5 6 100
R5 6 0 100
.OP
.ENDS
