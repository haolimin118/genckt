*scale(2)	circuit type(Clock RC tree (random fanout))

VIN 1 0 1
R0 1 2 100
C0 2 0 1p
R1 2 3 100
C1 3 0 1p
R2 2 4 100
C2 4 0 1p
R3 3 5 100
C3 5 0 1p
R4 4 6 100
C4 6 0 1p
R5 4 7 100
C5 7 0 1p
R6 5 8 100
C6 8 0 1p
R7 5 9 100
C7 9 0 1p
R8 6 10 100
C8 10 0 1p
R9 7 11 100
C9 11 0 1p
R10 7 12 100
C10 12 0 1p
R11 8 13 100
C11 13 0 1p
R12 8 14 100
C12 14 0 1p
R13 9 15 100
C13 15 0 1p
R14 10 16 100
C14 16 0 1p
R15 11 17 100
C15 17 0 1p
R16 12 18 100
C16 18 0 1p
R17 12 19 100
C17 19 0 1p
R18 13 20 100
C18 20 0 1p
R19 14 21 100
C19 21 0 1p
R20 15 22 100
C20 22 0 1p
R21 16 23 100
C21 23 0 1p
R22 17 24 100
C22 24 0 1p
R23 17 25 100
C23 25 0 1p
R24 18 26 100
C24 26 0 1p
R25 19 27 100
C25 27 0 1p
.OP
.ENDS
