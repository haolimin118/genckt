*scale(1)	circuit type(Mesh R)

VIN 1 0 1
R1 1 2 100
R2 1 3 100
R3 2 4 100
R4 3 4 100
R5 3 0 100

.OP
.PRINT V(3)
.ends
