*scale(2)	circuit type(Clock R tree (random fanout))

VIN 1 0 1
R0 1 2 100
R1 2 3 100
R2 2 4 100
R3 3 5 100
R4 3 6 100
R5 4 7 100
R6 5 8 100
R7 6 9 100
R8 6 10 100
R9 7 11 100
R10 7 12 100
R11 8 13 100
R12 9 14 100
R13 9 15 100
R14 10 16 100
R15 11 17 100
R16 12 18 100
R17 13 0 100
R18 13 0 100
R19 14 0 100
R20 15 0 100
R21 16 0 100
R22 17 0 100
R23 17 0 100
R24 18 0 100
R25 18 0 100
.OP
.ENDS
