*scale(50)	circuit type(RC ladder)

VIN 1 0 1
R1 1 2 100
C1 2 0 1p
R2 2 3 100
C2 3 0 1p
R3 3 4 100
C3 4 0 1p
R4 4 5 100
C4 5 0 1p
R5 5 6 100
C5 6 0 1p
R6 6 7 100
C6 7 0 1p
R7 7 8 100
C7 8 0 1p
R8 8 9 100
C8 9 0 1p
R9 9 10 100
C9 10 0 1p
R10 10 11 100
C10 11 0 1p
R11 11 12 100
C11 12 0 1p
R12 12 13 100
C12 13 0 1p
R13 13 14 100
C13 14 0 1p
R14 14 15 100
C14 15 0 1p
R15 15 16 100
C15 16 0 1p
R16 16 17 100
C16 17 0 1p
R17 17 18 100
C17 18 0 1p
R18 18 19 100
C18 19 0 1p
R19 19 20 100
C19 20 0 1p
R20 20 21 100
C20 21 0 1p
R21 21 22 100
C21 22 0 1p
R22 22 23 100
C22 23 0 1p
R23 23 24 100
C23 24 0 1p
R24 24 25 100
C24 25 0 1p
R25 25 26 100
C25 26 0 1p
R26 26 27 100
C26 27 0 1p
R27 27 28 100
C27 28 0 1p
R28 28 29 100
C28 29 0 1p
R29 29 30 100
C29 30 0 1p
R30 30 31 100
C30 31 0 1p
R31 31 32 100
C31 32 0 1p
R32 32 33 100
C32 33 0 1p
R33 33 34 100
C33 34 0 1p
R34 34 35 100
C34 35 0 1p
R35 35 36 100
C35 36 0 1p
R36 36 37 100
C36 37 0 1p
R37 37 38 100
C37 38 0 1p
R38 38 39 100
C38 39 0 1p
R39 39 40 100
C39 40 0 1p
R40 40 41 100
C40 41 0 1p
R41 41 42 100
C41 42 0 1p
R42 42 43 100
C42 43 0 1p
R43 43 44 100
C43 44 0 1p
R44 44 45 100
C44 45 0 1p
R45 45 46 100
C45 46 0 1p
R46 46 47 100
C46 47 0 1p
R47 47 48 100
C47 48 0 1p
R48 48 49 100
C48 49 0 1p
R49 49 50 100
C49 50 0 1p
R50 50 51 100
C50 51 0 1p

.OP
.PRINT V(51)
.ends
