*scale(5)	circuit type(Mesh R)

VIN 1 0 1
R1 1 2 100
R2 2 3 100
R3 3 4 100
R4 4 5 100
R5 5 6 100
R6 1 7 100
R7 2 8 100
R8 3 9 100
R9 4 10 100
R10 5 11 100
R11 6 12 100
R12 7 8 100
R13 8 9 100
R14 9 10 100
R15 10 11 100
R16 11 12 100
R17 7 13 100
R18 8 14 100
R19 9 15 100
R20 10 16 100
R21 11 17 100
R22 12 18 100
R23 13 14 100
R24 14 15 100
R25 15 16 100
R26 16 17 100
R27 17 18 100
R28 13 19 100
R29 14 20 100
R30 15 21 100
R31 16 22 100
R32 17 23 100
R33 18 24 100
R34 19 20 100
R35 20 21 100
R36 21 22 100
R37 22 23 100
R38 23 24 100
R39 19 25 100
R40 20 26 100
R41 21 27 100
R42 22 28 100
R43 23 29 100
R44 24 30 100
R45 25 26 100
R46 26 27 100
R47 27 28 100
R48 28 29 100
R49 29 30 100
R50 25 31 100
R51 26 32 100
R52 27 33 100
R53 28 34 100
R54 29 35 100
R55 30 36 100
R56 31 32 100
R57 32 33 100
R58 33 34 100
R59 34 35 100
R60 35 36 100
R61 31 0 100

.OP
.PRINT V(31)
.ends
