*scale (1), circuit type (ladderrc)

RC ladder --scale=1
VIN 1 0 1
R0 0 1 100
C0 1 0 1p
R1 1 2 100
C1 2 0 1p

.OP
.PRINT V(2)
.ends
