*scale(2)	circuit type(Mesh R)

VIN 1 0 1
R1 1 2 100
R2 2 3 100
R3 1 4 100
R4 2 5 100
R5 3 6 100
R6 4 5 100
R7 5 6 100
R8 4 7 100
R9 5 8 100
R10 6 9 100
R11 7 8 100
R12 8 9 100
R13 7 0 100

.OP
.PRINT V(7)
.ends
