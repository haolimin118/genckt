*scale (5), circuit type (ladderrlc)

RLC ladder --scale=5
VIN 1 0 1
C0 1 0 1p
R1 1 2 100
L1 2 3 1m
C1 3 0 1p
R2 3 4 100
L2 4 5 1m
C2 5 0 1p
R3 5 6 100
L3 6 7 1m
C3 7 0 1p
R4 7 8 100
L4 8 9 1m
C4 9 0 1p
R5 9 10 100
L5 10 11 1m
C5 11 0 1p

.OP
.PRINT V(11)
.ends
