*scale (1), circuit type (ladderrc)

VIN 1 0 1
R1 1 2 100
C1 2 0 1p

.OP
.PRINT V(2)
.ends
