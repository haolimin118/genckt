*scale(2)	circuit type(Clock R tree)

VIN 1 0 1
R0 1 2 100
R1 2 3 100
R2 2 4 100
R3 3 5 100
R4 3 6 100
R5 4 7 100
R6 4 8 100
R7 5 9 100
R8 5 10 100
R9 6 11 100
R10 6 12 100
R11 7 13 100
R12 7 14 100
R13 8 15 100
R14 8 16 100
R15 9 17 100
R16 9 18 100
R17 10 19 100
R18 10 20 100
R19 11 21 100
R20 11 22 100
R21 12 23 100
R22 12 24 100
R23 13 25 100
R24 13 26 100
R25 14 27 100
R26 14 28 100
R27 15 29 100
R28 15 30 100
R29 16 31 100
R30 16 32 100
R31 17 0 100
R32 17 0 100
R33 18 0 100
R34 18 0 100
R35 19 0 100
R36 19 0 100
R37 20 0 100
R38 20 0 100
R39 21 0 100
R40 21 0 100
R41 22 0 100
R42 22 0 100
R43 23 0 100
R44 23 0 100
R45 24 0 100
R46 24 0 100
R47 25 0 100
R48 25 0 100
R49 26 0 100
R50 26 0 100
R51 27 0 100
R52 27 0 100
R53 28 0 100
R54 28 0 100
R55 29 0 100
R56 29 0 100
R57 30 0 100
R58 30 0 100
R59 31 0 100
R60 31 0 100
R61 32 0 100
R62 32 0 100
.OP
.ENDS
